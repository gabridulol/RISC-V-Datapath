`include "PC.v"

module Datapath (
    input wire clock, reset,


);

endmodule

module Datapath_Testbench;



endmodule