module Datapath (

)

endmodule